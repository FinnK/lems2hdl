izhikevichCell-