iafRefCell-