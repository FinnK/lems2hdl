pointCellCondBased-channelPopulation-ionChannelPassive-channelPopulation-ionChannelHH-gateHHrates-HHExpLinearRate-HHExpRate-gateHHrates-HHExpRate-HHSigmoidRate-channelPopulation-ionChannelHH-gateHHrates-HHExpLinearRate-HHExpRate-